/*
 * Copyright (c) 2025 Toivo Henningsson
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module pulse_width_modulator #(
		parameter BITS=11
	) (
		input wire clk, reset,

		input wire dual_slope_en, double_slope_en, ddr_en,
		input wire [BITS-1:0] compare_max, // controls the PWM period, pulse_width should be <= compare_max (less if´one pulse/period is wanted)

		input wire [BITS-1:0] pulse_width, // range is -1/4*2^BITS <= pulse_width < 3/4*2^BITS
		output wire pulse_done, // when high, supply the next pulse_width value in the next cycle
		output wire pwm_out
	);

	reg direction;
	reg [BITS-1:0] compare_value;

	//wire compare_value_at_max = (compare_value == compare_max);
	// To avoid taking a very long period when changing compare value. We could reset the compare value instead when changing compare_max?
	wire compare_value_at_max = compare_value >= compare_max;

	// not registers
	reg r_restart, r_pulse_done;
	reg signed [2:0] delta;
	reg next_direction;
	always_comb begin
		if (dual_slope_en) begin
			delta = direction ? 1 : -1;
			if (double_slope_en) delta = direction ? 2 : -2;

			next_direction = direction;
			if (compare_value_at_max && (direction == 1)) begin
				delta = double_slope_en ? -1 : 0;
				next_direction = 0;
			end

			r_restart = (direction == 0) && (compare_value[BITS-1:1] == 0) && (double_slope_en || compare_value[0] == 0);
			r_pulse_done = (direction == 1) && compare_value_at_max;
		end else begin
			delta = double_slope_en ? 2 : 1;
			next_direction = 1;

			r_restart = compare_value_at_max;
			r_pulse_done = r_restart;
		end
	end
//	assign pulse_done = r_restart;
	assign pulse_done = r_pulse_done;

	always_ff @(posedge clk) begin
		if (reset) begin
			direction <= 1;
			compare_value <= double_slope_en;
		end else begin
			if (r_restart) compare_value <= double_slope_en;
			else compare_value <= $signed(compare_value) + $signed(delta);

			direction <= r_restart ? 1 : next_direction;
		end
	end

	// TODO: Hold the pulse together? Now it's the low pulse that is continuous -- shouldn't make a difference though
	//assign pwm_out = pulse_width[BITS-1] ? !pulse_width[BITS-2] : (compare_value < pulse_width);

	wire pwm_cmp = (compare_value < pulse_width);
	wire pwm_eq = (compare_value == pulse_width);

	wire pwm1_0 = pwm_cmp || (ddr_en && pwm_eq && pulse_width[0]);
	wire pwm2_0 = pwm_cmp || (ddr_en && pwm_eq && !pulse_width[0]);

	wire pwm1 = pulse_width[BITS-1] ? !pulse_width[BITS-2] : pwm1_0;
	wire pwm2 = pulse_width[BITS-1] ? !pulse_width[BITS-2] : pwm2_0;

	/*
	reg pwm_reg;
	always_ff @(posedge clk) pwm_reg <= pwm1;
	assign pwm_out = pwm_reg;
	*/
	
	reg pwm_reg, pwm_reg_n;
	always_ff @(posedge clk) pwm_reg <= !pwm2;

	//always_ff @(negedge clk) pwm_reg_n <= !pwm1 | !ddr_en; // Note: negedge
	//assign pwm_out = !(pwm_reg & pwm_reg_n);

	always_ff @(negedge clk) pwm_reg_n <= !pwm1 && ddr_en; // Note: negedge
	assign pwm_out = !(pwm_reg || pwm_reg_n);
endmodule : pulse_width_modulator
